module verilog_practice (input A , B, output S, C);
//Structure Modelling
xor(S,A,B);
and(C,A,B);
///

// Data dlow modeling
//assign S = A^B;
//assign C= A&B;

//

endmodule 